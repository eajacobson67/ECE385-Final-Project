typedef logic [2:0] [31:0] vector;
typedef logic [31:0] fixed_real;
typedef logic [2:0] [31:0] color;

module y_ang_lut (
	input logic Clk,
	input logic [9:0] WriteY,
	output fixed_real dPhi
);

logic [9:0] in_0;
logic [8:0] in;
logic [15:0] out, out_signed;

assign in_0 = (WriteY >= 10'd240)?WriteY-10'd240:10'd240-WriteY;
assign in = in_0[8:0];
assign out_signed = (WriteY >= 10'd240)?out:(~out)+1;
assign dPhi = {out_signed,16'b0};

/*
function tobin(a){
	var str = Math.round(a);
	return str.toString(2);
}

var out = "always_ff @ (negedge Clk) begin\ncase (in)\n";
for(var i = 0; i <= 240; i++) {
		out += "9'd" + (i) + ": out <= 16'b"+tobin(Math.atan(i/240)/Math.PI*180)+";    ";
		if(!(i % 3)){
			out += "\n";
		}
}
out += "endcase\nend\n";
console.log(out);
*/
always_ff @ (negedge Clk) begin
case (in)
9'd0: out <= 16'b0;    
9'd1: out <= 16'b0;    9'd2: out <= 16'b0;    9'd3: out <= 16'b1;    
9'd4: out <= 16'b1;    9'd5: out <= 16'b1;    9'd6: out <= 16'b1;    
9'd7: out <= 16'b10;    9'd8: out <= 16'b10;    9'd9: out <= 16'b10;    
9'd10: out <= 16'b10;    9'd11: out <= 16'b11;    9'd12: out <= 16'b11;    
9'd13: out <= 16'b11;    9'd14: out <= 16'b11;    9'd15: out <= 16'b100;    
9'd16: out <= 16'b100;    9'd17: out <= 16'b100;    9'd18: out <= 16'b100;    
9'd19: out <= 16'b101;    9'd20: out <= 16'b101;    9'd21: out <= 16'b101;    
9'd22: out <= 16'b101;    9'd23: out <= 16'b101;    9'd24: out <= 16'b110;    
9'd25: out <= 16'b110;    9'd26: out <= 16'b110;    9'd27: out <= 16'b110;    
9'd28: out <= 16'b111;    9'd29: out <= 16'b111;    9'd30: out <= 16'b111;    
9'd31: out <= 16'b111;    9'd32: out <= 16'b1000;    9'd33: out <= 16'b1000;    
9'd34: out <= 16'b1000;    9'd35: out <= 16'b1000;    9'd36: out <= 16'b1001;    
9'd37: out <= 16'b1001;    9'd38: out <= 16'b1001;    9'd39: out <= 16'b1001;    
9'd40: out <= 16'b1001;    9'd41: out <= 16'b1010;    9'd42: out <= 16'b1010;    
9'd43: out <= 16'b1010;    9'd44: out <= 16'b1010;    9'd45: out <= 16'b1011;    
9'd46: out <= 16'b1011;    9'd47: out <= 16'b1011;    9'd48: out <= 16'b1011;    
9'd49: out <= 16'b1100;    9'd50: out <= 16'b1100;    9'd51: out <= 16'b1100;    
9'd52: out <= 16'b1100;    9'd53: out <= 16'b1100;    9'd54: out <= 16'b1101;    
9'd55: out <= 16'b1101;    9'd56: out <= 16'b1101;    9'd57: out <= 16'b1101;    
9'd58: out <= 16'b1110;    9'd59: out <= 16'b1110;    9'd60: out <= 16'b1110;    
9'd61: out <= 16'b1110;    9'd62: out <= 16'b1110;    9'd63: out <= 16'b1111;    
9'd64: out <= 16'b1111;    9'd65: out <= 16'b1111;    9'd66: out <= 16'b1111;    
9'd67: out <= 16'b10000;    9'd68: out <= 16'b10000;    9'd69: out <= 16'b10000;    
9'd70: out <= 16'b10000;    9'd71: out <= 16'b10000;    9'd72: out <= 16'b10001;    
9'd73: out <= 16'b10001;    9'd74: out <= 16'b10001;    9'd75: out <= 16'b10001;    
9'd76: out <= 16'b10010;    9'd77: out <= 16'b10010;    9'd78: out <= 16'b10010;    
9'd79: out <= 16'b10010;    9'd80: out <= 16'b10010;    9'd81: out <= 16'b10011;    
9'd82: out <= 16'b10011;    9'd83: out <= 16'b10011;    9'd84: out <= 16'b10011;    
9'd85: out <= 16'b10100;    9'd86: out <= 16'b10100;    9'd87: out <= 16'b10100;    
9'd88: out <= 16'b10100;    9'd89: out <= 16'b10100;    9'd90: out <= 16'b10101;    
9'd91: out <= 16'b10101;    9'd92: out <= 16'b10101;    9'd93: out <= 16'b10101;    
9'd94: out <= 16'b10101;    9'd95: out <= 16'b10110;    9'd96: out <= 16'b10110;    
9'd97: out <= 16'b10110;    9'd98: out <= 16'b10110;    9'd99: out <= 16'b10110;    
9'd100: out <= 16'b10111;    9'd101: out <= 16'b10111;    9'd102: out <= 16'b10111;    
9'd103: out <= 16'b10111;    9'd104: out <= 16'b10111;    9'd105: out <= 16'b11000;    
9'd106: out <= 16'b11000;    9'd107: out <= 16'b11000;    9'd108: out <= 16'b11000;    
9'd109: out <= 16'b11000;    9'd110: out <= 16'b11001;    9'd111: out <= 16'b11001;    
9'd112: out <= 16'b11001;    9'd113: out <= 16'b11001;    9'd114: out <= 16'b11001;    
9'd115: out <= 16'b11010;    9'd116: out <= 16'b11010;    9'd117: out <= 16'b11010;    
9'd118: out <= 16'b11010;    9'd119: out <= 16'b11010;    9'd120: out <= 16'b11011;    
9'd121: out <= 16'b11011;    9'd122: out <= 16'b11011;    9'd123: out <= 16'b11011;    
9'd124: out <= 16'b11011;    9'd125: out <= 16'b11100;    9'd126: out <= 16'b11100;    
9'd127: out <= 16'b11100;    9'd128: out <= 16'b11100;    9'd129: out <= 16'b11100;    
9'd130: out <= 16'b11100;    9'd131: out <= 16'b11101;    9'd132: out <= 16'b11101;    
9'd133: out <= 16'b11101;    9'd134: out <= 16'b11101;    9'd135: out <= 16'b11101;    
9'd136: out <= 16'b11110;    9'd137: out <= 16'b11110;    9'd138: out <= 16'b11110;    
9'd139: out <= 16'b11110;    9'd140: out <= 16'b11110;    9'd141: out <= 16'b11110;    
9'd142: out <= 16'b11111;    9'd143: out <= 16'b11111;    9'd144: out <= 16'b11111;    
9'd145: out <= 16'b11111;    9'd146: out <= 16'b11111;    9'd147: out <= 16'b11111;    
9'd148: out <= 16'b100000;    9'd149: out <= 16'b100000;    9'd150: out <= 16'b100000;    
9'd151: out <= 16'b100000;    9'd152: out <= 16'b100000;    9'd153: out <= 16'b100001;    
9'd154: out <= 16'b100001;    9'd155: out <= 16'b100001;    9'd156: out <= 16'b100001;    
9'd157: out <= 16'b100001;    9'd158: out <= 16'b100001;    9'd159: out <= 16'b100010;    
9'd160: out <= 16'b100010;    9'd161: out <= 16'b100010;    9'd162: out <= 16'b100010;    
9'd163: out <= 16'b100010;    9'd164: out <= 16'b100010;    9'd165: out <= 16'b100011;    
9'd166: out <= 16'b100011;    9'd167: out <= 16'b100011;    9'd168: out <= 16'b100011;    
9'd169: out <= 16'b100011;    9'd170: out <= 16'b100011;    9'd171: out <= 16'b100011;    
9'd172: out <= 16'b100100;    9'd173: out <= 16'b100100;    9'd174: out <= 16'b100100;    
9'd175: out <= 16'b100100;    9'd176: out <= 16'b100100;    9'd177: out <= 16'b100100;    
9'd178: out <= 16'b100101;    9'd179: out <= 16'b100101;    9'd180: out <= 16'b100101;    
9'd181: out <= 16'b100101;    9'd182: out <= 16'b100101;    9'd183: out <= 16'b100101;    
9'd184: out <= 16'b100101;    9'd185: out <= 16'b100110;    9'd186: out <= 16'b100110;    
9'd187: out <= 16'b100110;    9'd188: out <= 16'b100110;    9'd189: out <= 16'b100110;    
9'd190: out <= 16'b100110;    9'd191: out <= 16'b100111;    9'd192: out <= 16'b100111;    
9'd193: out <= 16'b100111;    9'd194: out <= 16'b100111;    9'd195: out <= 16'b100111;    
9'd196: out <= 16'b100111;    9'd197: out <= 16'b100111;    9'd198: out <= 16'b101000;    
9'd199: out <= 16'b101000;    9'd200: out <= 16'b101000;    9'd201: out <= 16'b101000;    
9'd202: out <= 16'b101000;    9'd203: out <= 16'b101000;    9'd204: out <= 16'b101000;    
9'd205: out <= 16'b101001;    9'd206: out <= 16'b101001;    9'd207: out <= 16'b101001;    
9'd208: out <= 16'b101001;    9'd209: out <= 16'b101001;    9'd210: out <= 16'b101001;    
9'd211: out <= 16'b101001;    9'd212: out <= 16'b101001;    9'd213: out <= 16'b101010;    
9'd214: out <= 16'b101010;    9'd215: out <= 16'b101010;    9'd216: out <= 16'b101010;    
9'd217: out <= 16'b101010;    9'd218: out <= 16'b101010;    9'd219: out <= 16'b101010;    
9'd220: out <= 16'b101011;    9'd221: out <= 16'b101011;    9'd222: out <= 16'b101011;    
9'd223: out <= 16'b101011;    9'd224: out <= 16'b101011;    9'd225: out <= 16'b101011;    
9'd226: out <= 16'b101011;    9'd227: out <= 16'b101011;    9'd228: out <= 16'b101100;    
9'd229: out <= 16'b101100;    9'd230: out <= 16'b101100;    9'd231: out <= 16'b101100;    
9'd232: out <= 16'b101100;    9'd233: out <= 16'b101100;    9'd234: out <= 16'b101100;    
9'd235: out <= 16'b101100;    9'd236: out <= 16'b101101;    9'd237: out <= 16'b101101;    
9'd238: out <= 16'b101101;    9'd239: out <= 16'b101101;    9'd240: out <= 16'b101101;    
endcase

end


endmodule

module x_ang_lut (
	input logic Clk,
	input logic [9:0] WriteX,
	output fixed_real dTheta
);

logic [9:0] in_0;
logic [8:0] in;
logic [15:0] out, out_signed;

assign in_0 = (WriteX >= 10'd320)?WriteX-10'd320:10'd320-WriteX;
assign in = in_0[8:0];
assign out_signed = (WriteX > 10'd320)?(~out)+1:out;
assign dTheta = {out_signed,16'b0};

/*
function tobin(a){
	var str = Math.round(a);
	return str.toString(2);
}

var out = "always_ff @ (negedge Clk) begin\ncase (in)\n";
for(var i = 0; i <= 320; i++) {
		out += "9'd" + (i) + ": out <= 16'b"+tobin(Math.atan(i/240)/Math.PI*180)+";    ";
		if(!(i % 3)){
			out += "\n";
		}
}
out += "endcase\nend\n";
console.log(out);
*/
always_ff @ (negedge Clk) begin
case (in)
9'd0: out <= 16'b0;    
9'd1: out <= 16'b0;    9'd2: out <= 16'b0;    9'd3: out <= 16'b1;    
9'd4: out <= 16'b1;    9'd5: out <= 16'b1;    9'd6: out <= 16'b1;    
9'd7: out <= 16'b10;    9'd8: out <= 16'b10;    9'd9: out <= 16'b10;    
9'd10: out <= 16'b10;    9'd11: out <= 16'b11;    9'd12: out <= 16'b11;    
9'd13: out <= 16'b11;    9'd14: out <= 16'b11;    9'd15: out <= 16'b100;    
9'd16: out <= 16'b100;    9'd17: out <= 16'b100;    9'd18: out <= 16'b100;    
9'd19: out <= 16'b101;    9'd20: out <= 16'b101;    9'd21: out <= 16'b101;    
9'd22: out <= 16'b101;    9'd23: out <= 16'b101;    9'd24: out <= 16'b110;    
9'd25: out <= 16'b110;    9'd26: out <= 16'b110;    9'd27: out <= 16'b110;    
9'd28: out <= 16'b111;    9'd29: out <= 16'b111;    9'd30: out <= 16'b111;    
9'd31: out <= 16'b111;    9'd32: out <= 16'b1000;    9'd33: out <= 16'b1000;    
9'd34: out <= 16'b1000;    9'd35: out <= 16'b1000;    9'd36: out <= 16'b1001;    
9'd37: out <= 16'b1001;    9'd38: out <= 16'b1001;    9'd39: out <= 16'b1001;    
9'd40: out <= 16'b1001;    9'd41: out <= 16'b1010;    9'd42: out <= 16'b1010;    
9'd43: out <= 16'b1010;    9'd44: out <= 16'b1010;    9'd45: out <= 16'b1011;    
9'd46: out <= 16'b1011;    9'd47: out <= 16'b1011;    9'd48: out <= 16'b1011;    
9'd49: out <= 16'b1100;    9'd50: out <= 16'b1100;    9'd51: out <= 16'b1100;    
9'd52: out <= 16'b1100;    9'd53: out <= 16'b1100;    9'd54: out <= 16'b1101;    
9'd55: out <= 16'b1101;    9'd56: out <= 16'b1101;    9'd57: out <= 16'b1101;    
9'd58: out <= 16'b1110;    9'd59: out <= 16'b1110;    9'd60: out <= 16'b1110;    
9'd61: out <= 16'b1110;    9'd62: out <= 16'b1110;    9'd63: out <= 16'b1111;    
9'd64: out <= 16'b1111;    9'd65: out <= 16'b1111;    9'd66: out <= 16'b1111;    
9'd67: out <= 16'b10000;    9'd68: out <= 16'b10000;    9'd69: out <= 16'b10000;    
9'd70: out <= 16'b10000;    9'd71: out <= 16'b10000;    9'd72: out <= 16'b10001;    
9'd73: out <= 16'b10001;    9'd74: out <= 16'b10001;    9'd75: out <= 16'b10001;    
9'd76: out <= 16'b10010;    9'd77: out <= 16'b10010;    9'd78: out <= 16'b10010;    
9'd79: out <= 16'b10010;    9'd80: out <= 16'b10010;    9'd81: out <= 16'b10011;    
9'd82: out <= 16'b10011;    9'd83: out <= 16'b10011;    9'd84: out <= 16'b10011;    
9'd85: out <= 16'b10100;    9'd86: out <= 16'b10100;    9'd87: out <= 16'b10100;    
9'd88: out <= 16'b10100;    9'd89: out <= 16'b10100;    9'd90: out <= 16'b10101;    
9'd91: out <= 16'b10101;    9'd92: out <= 16'b10101;    9'd93: out <= 16'b10101;    
9'd94: out <= 16'b10101;    9'd95: out <= 16'b10110;    9'd96: out <= 16'b10110;    
9'd97: out <= 16'b10110;    9'd98: out <= 16'b10110;    9'd99: out <= 16'b10110;    
9'd100: out <= 16'b10111;    9'd101: out <= 16'b10111;    9'd102: out <= 16'b10111;    
9'd103: out <= 16'b10111;    9'd104: out <= 16'b10111;    9'd105: out <= 16'b11000;    
9'd106: out <= 16'b11000;    9'd107: out <= 16'b11000;    9'd108: out <= 16'b11000;    
9'd109: out <= 16'b11000;    9'd110: out <= 16'b11001;    9'd111: out <= 16'b11001;    
9'd112: out <= 16'b11001;    9'd113: out <= 16'b11001;    9'd114: out <= 16'b11001;    
9'd115: out <= 16'b11010;    9'd116: out <= 16'b11010;    9'd117: out <= 16'b11010;    
9'd118: out <= 16'b11010;    9'd119: out <= 16'b11010;    9'd120: out <= 16'b11011;    
9'd121: out <= 16'b11011;    9'd122: out <= 16'b11011;    9'd123: out <= 16'b11011;    
9'd124: out <= 16'b11011;    9'd125: out <= 16'b11100;    9'd126: out <= 16'b11100;    
9'd127: out <= 16'b11100;    9'd128: out <= 16'b11100;    9'd129: out <= 16'b11100;    
9'd130: out <= 16'b11100;    9'd131: out <= 16'b11101;    9'd132: out <= 16'b11101;    
9'd133: out <= 16'b11101;    9'd134: out <= 16'b11101;    9'd135: out <= 16'b11101;    
9'd136: out <= 16'b11110;    9'd137: out <= 16'b11110;    9'd138: out <= 16'b11110;    
9'd139: out <= 16'b11110;    9'd140: out <= 16'b11110;    9'd141: out <= 16'b11110;    
9'd142: out <= 16'b11111;    9'd143: out <= 16'b11111;    9'd144: out <= 16'b11111;    
9'd145: out <= 16'b11111;    9'd146: out <= 16'b11111;    9'd147: out <= 16'b11111;    
9'd148: out <= 16'b100000;    9'd149: out <= 16'b100000;    9'd150: out <= 16'b100000;    
9'd151: out <= 16'b100000;    9'd152: out <= 16'b100000;    9'd153: out <= 16'b100001;    
9'd154: out <= 16'b100001;    9'd155: out <= 16'b100001;    9'd156: out <= 16'b100001;    
9'd157: out <= 16'b100001;    9'd158: out <= 16'b100001;    9'd159: out <= 16'b100010;    
9'd160: out <= 16'b100010;    9'd161: out <= 16'b100010;    9'd162: out <= 16'b100010;    
9'd163: out <= 16'b100010;    9'd164: out <= 16'b100010;    9'd165: out <= 16'b100011;    
9'd166: out <= 16'b100011;    9'd167: out <= 16'b100011;    9'd168: out <= 16'b100011;    
9'd169: out <= 16'b100011;    9'd170: out <= 16'b100011;    9'd171: out <= 16'b100011;    
9'd172: out <= 16'b100100;    9'd173: out <= 16'b100100;    9'd174: out <= 16'b100100;    
9'd175: out <= 16'b100100;    9'd176: out <= 16'b100100;    9'd177: out <= 16'b100100;    
9'd178: out <= 16'b100101;    9'd179: out <= 16'b100101;    9'd180: out <= 16'b100101;    
9'd181: out <= 16'b100101;    9'd182: out <= 16'b100101;    9'd183: out <= 16'b100101;    
9'd184: out <= 16'b100101;    9'd185: out <= 16'b100110;    9'd186: out <= 16'b100110;    
9'd187: out <= 16'b100110;    9'd188: out <= 16'b100110;    9'd189: out <= 16'b100110;    
9'd190: out <= 16'b100110;    9'd191: out <= 16'b100111;    9'd192: out <= 16'b100111;    
9'd193: out <= 16'b100111;    9'd194: out <= 16'b100111;    9'd195: out <= 16'b100111;    
9'd196: out <= 16'b100111;    9'd197: out <= 16'b100111;    9'd198: out <= 16'b101000;    
9'd199: out <= 16'b101000;    9'd200: out <= 16'b101000;    9'd201: out <= 16'b101000;    
9'd202: out <= 16'b101000;    9'd203: out <= 16'b101000;    9'd204: out <= 16'b101000;    
9'd205: out <= 16'b101001;    9'd206: out <= 16'b101001;    9'd207: out <= 16'b101001;    
9'd208: out <= 16'b101001;    9'd209: out <= 16'b101001;    9'd210: out <= 16'b101001;    
9'd211: out <= 16'b101001;    9'd212: out <= 16'b101001;    9'd213: out <= 16'b101010;    
9'd214: out <= 16'b101010;    9'd215: out <= 16'b101010;    9'd216: out <= 16'b101010;    
9'd217: out <= 16'b101010;    9'd218: out <= 16'b101010;    9'd219: out <= 16'b101010;    
9'd220: out <= 16'b101011;    9'd221: out <= 16'b101011;    9'd222: out <= 16'b101011;    
9'd223: out <= 16'b101011;    9'd224: out <= 16'b101011;    9'd225: out <= 16'b101011;    
9'd226: out <= 16'b101011;    9'd227: out <= 16'b101011;    9'd228: out <= 16'b101100;    
9'd229: out <= 16'b101100;    9'd230: out <= 16'b101100;    9'd231: out <= 16'b101100;    
9'd232: out <= 16'b101100;    9'd233: out <= 16'b101100;    9'd234: out <= 16'b101100;    
9'd235: out <= 16'b101100;    9'd236: out <= 16'b101101;    9'd237: out <= 16'b101101;    
9'd238: out <= 16'b101101;    9'd239: out <= 16'b101101;    9'd240: out <= 16'b101101;    
9'd241: out <= 16'b101101;    9'd242: out <= 16'b101101;    9'd243: out <= 16'b101101;    
9'd244: out <= 16'b101101;    9'd245: out <= 16'b101110;    9'd246: out <= 16'b101110;    
9'd247: out <= 16'b101110;    9'd248: out <= 16'b101110;    9'd249: out <= 16'b101110;    
9'd250: out <= 16'b101110;    9'd251: out <= 16'b101110;    9'd252: out <= 16'b101110;    
9'd253: out <= 16'b101111;    9'd254: out <= 16'b101111;    9'd255: out <= 16'b101111;    
9'd256: out <= 16'b101111;    9'd257: out <= 16'b101111;    9'd258: out <= 16'b101111;    
9'd259: out <= 16'b101111;    9'd260: out <= 16'b101111;    9'd261: out <= 16'b101111;    
9'd262: out <= 16'b110000;    9'd263: out <= 16'b110000;    9'd264: out <= 16'b110000;    
9'd265: out <= 16'b110000;    9'd266: out <= 16'b110000;    9'd267: out <= 16'b110000;    
9'd268: out <= 16'b110000;    9'd269: out <= 16'b110000;    9'd270: out <= 16'b110000;    
9'd271: out <= 16'b110000;    9'd272: out <= 16'b110001;    9'd273: out <= 16'b110001;    
9'd274: out <= 16'b110001;    9'd275: out <= 16'b110001;    9'd276: out <= 16'b110001;    
9'd277: out <= 16'b110001;    9'd278: out <= 16'b110001;    9'd279: out <= 16'b110001;    
9'd280: out <= 16'b110001;    9'd281: out <= 16'b110001;    9'd282: out <= 16'b110010;    
9'd283: out <= 16'b110010;    9'd284: out <= 16'b110010;    9'd285: out <= 16'b110010;    
9'd286: out <= 16'b110010;    9'd287: out <= 16'b110010;    9'd288: out <= 16'b110010;    
9'd289: out <= 16'b110010;    9'd290: out <= 16'b110010;    9'd291: out <= 16'b110010;    
9'd292: out <= 16'b110011;    9'd293: out <= 16'b110011;    9'd294: out <= 16'b110011;    
9'd295: out <= 16'b110011;    9'd296: out <= 16'b110011;    9'd297: out <= 16'b110011;    
9'd298: out <= 16'b110011;    9'd299: out <= 16'b110011;    9'd300: out <= 16'b110011;    
9'd301: out <= 16'b110011;    9'd302: out <= 16'b110100;    9'd303: out <= 16'b110100;    
9'd304: out <= 16'b110100;    9'd305: out <= 16'b110100;    9'd306: out <= 16'b110100;    
9'd307: out <= 16'b110100;    9'd308: out <= 16'b110100;    9'd309: out <= 16'b110100;    
9'd310: out <= 16'b110100;    9'd311: out <= 16'b110100;    9'd312: out <= 16'b110100;    
9'd313: out <= 16'b110101;    9'd314: out <= 16'b110101;    9'd315: out <= 16'b110101;    
9'd316: out <= 16'b110101;    9'd317: out <= 16'b110101;    9'd318: out <= 16'b110101;    
9'd319: out <= 16'b110101;    9'd320: out <= 16'b110101;    endcase
end

endmodule
